------------------------------------------------------------------------------
--  LEON3 Demonstration design
--  Copyright (C) 2006 Jiri Gaisler, Gaisler Research
------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2014, Aeroflex Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library grlib;
use grlib.config.all;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;
library techmap;
use techmap.gencomp.all;
use techmap.allclkgen.all;
library gaisler;
use gaisler.memctrl.all;
use gaisler.leon3.all;
use gaisler.uart.all;
use gaisler.misc.all;
use gaisler.i2c.all;
use gaisler.net.all;
use gaisler.jtag.all;
library esa;
use esa.memoryctrl.all;
use work.config.all;
use work.ml605.all;
-- pragma translate_off
use gaisler.sim.all;
-- pragma translate_on
library rvex;
use rvex.common_pkg.all;
use rvex.bus_pkg.all;
use rvex.bus_addrConv_pkg.all;
use rvex.core_pkg.all;
use rvex.cache_pkg.all;
use rvex.rvsys_grlib_pkg.all;
-- pragma translate_off
use rvex.utils_pkg.all;
use rvex.simUtils_pkg.all;
use rvex.simUtils_mem_pkg.all;
-- pragma translate_on
library unisim;
use unisim.vcomponents.all;
library work;
use work.platform_version_pkg.all;

entity leon3mp is
  generic (
    fabtech  : integer := CFG_FABTECH;
    memtech  : integer := CFG_MEMTECH;
    padtech  : integer := CFG_PADTECH;
    SIM_BYPASS_INIT_CAL : string := "OFF";
    DISABLE_DDR_SIM : boolean := false
  );
  port (
    
    -- System control.
    reset                       : in    std_ulogic;
    clk_ref_p                   : in    std_logic; -- 200 MHz.
    clk_ref_n                   : in    std_logic;
    gmiiclk_p                   : in    std_ulogic; -- 125 MHz.
    gmiiclk_n                   : in    std_ulogic;
    clk_33                      : in    std_ulogic; -- 33 MHz.
    
    -- DDR3 memory.
    ddr3_dq                     : inout std_logic_vector(DQ_WIDTH-1 downto 0);
    ddr3_dm                     : out   std_logic_vector(DM_WIDTH-1 downto 0);
    ddr3_addr                   : out   std_logic_vector(ROW_WIDTH-1 downto 0);
    ddr3_ba                     : out   std_logic_vector(BANK_WIDTH-1 downto 0);
    ddr3_ras_n                  : out   std_logic;
    ddr3_cas_n                  : out   std_logic;
    ddr3_we_n                   : out   std_logic;
    ddr3_reset_n                : out   std_logic;
    ddr3_cs_n                   : out   std_logic_vector((CS_WIDTH*nCS_PER_RANK)-1 downto 0);
    ddr3_odt                    : out   std_logic_vector((CS_WIDTH*nCS_PER_RANK)-1 downto 0);
    ddr3_cke                    : out   std_logic_vector(CKE_WIDTH-1 downto 0);
    ddr3_dqs_p                  : inout std_logic_vector(DQS_WIDTH-1 downto 0);
    ddr3_dqs_n                  : inout std_logic_vector(DQS_WIDTH-1 downto 0);
    ddr3_ck_p                   : out   std_logic_vector(CK_WIDTH-1 downto 0);
    ddr3_ck_n                   : out   std_logic_vector(CK_WIDTH-1 downto 0);

    -- Debug UART.
    dsurx                       : in    std_ulogic;
    dsutx                       : out   std_ulogic;
    
    -- GPIO.
    led                         : inout std_logic_vector(12 downto 0) := (others => '0'); -- LEDs (1..8, CWESN)
    dipsw                       : in    std_logic_vector(7 downto 0)  := (others => '0'); -- DIP switches (1..8)
    pbtn                        : in    std_logic_vector(4 downto 0)  := (others => '0')  -- Pushbuttons (CWESN)
    
  );
end;

architecture rtl of leon3mp is
  
  -- Attribute declarations.
  attribute keep                  : boolean;
  attribute syn_keep              : boolean;
  attribute syn_preserve          : boolean;
  
  -- Clocks.
  constant VCO_FREQ               : integer := 1200000; -- MMCM VCO frequency in KHz
  
  signal clk125                   : std_ulogic; -- 125 MHz from ethernet osc.
  signal clk100                   : std_ulogic; -- 100 MHz clock generated by the MIG.
  signal clk33                    : std_ulogic; -- 33 MHz from sysACE osc.
  
  signal clkm                     : std_ulogic;
  attribute syn_keep       of clkm: signal is true;
  attribute syn_preserve   of clkm: signal is true;
  attribute keep           of clkm: signal is true;
  constant CLKM_FREQ              : integer := VCO_FREQ / CFG_MIG_CLK4;
  
  -- PPL lock/reset bullshit.
  signal rstn                     : std_ulogic;
  signal rstraw                   : std_logic;
  signal lock                     : std_logic;
  attribute syn_keep       of lock: signal is true;
  attribute keep           of lock: signal is true;
  
  -- Memory controller stuff.
  signal migi		                  : mig_app_in_type;
  signal migo		                  : mig_app_out_type;
  signal clkddr                   : std_ulogic;
  attribute syn_keep     of clkddr: signal is true;
  attribute syn_preserve of clkddr: signal is true;
  attribute keep         of clkddr: signal is true;
  signal phy_init_done            : std_logic;

  -- AHB/APB/r-VEX bus.
  constant N_RVB_SLAVES           : integer := CFG_NRVEX + 3;
  signal apbi                     : apb_slv_in_type;
  signal apbo                     : apb_slv_out_vector := (others => apb_none);
  signal ahbsi                    : ahb_slv_in_type;
  signal ahbso                    : ahb_slv_out_vector := (others => ahbs_none);
  signal ahbmi                    : ahb_mst_in_type;
  signal ahbmo                    : ahb_mst_out_vector := (others => ahbm_none);
  signal rvbmo                    : bus_mst2slv_type;
  signal rvbmi                    : bus_slv2mst_type;
  signal rvbsi                    : bus_mst2slv_array(0 to N_RVB_SLAVES - 1);
  signal rvbso                    : bus_slv2mst_array(0 to N_RVB_SLAVES - 1);
  
  -- Interrupt requests.
  constant NIRQ                   : natural := 2;
  signal irq                      : std_logic_vector(NIRQ downto 1) := (others => '0');
  
  -- Interrupt control/r-VEX interface signals.
  signal irq2rv_irq               : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal irq2rv_irqID             : rvex_address_array(CFG_NCTXT-1 downto 0);
  signal rv2irq_irqAck            : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal busy2rv_run              : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal irq2busy_run             : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal rv2irq_idle              : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal rv2irq_break             : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal irq2rv_reset             : std_logic_vector(CFG_NCTXT-1 downto 0);
  signal irq2rv_resetVect         : rvex_address_array(CFG_NCTXT-1 downto 0);
  signal rv2irq_done              : std_logic_vector(CFG_NCTXT-1 downto 0);
  
  -- Trace stall broadcasting signals.
  signal rv2rctrl_traceStall      : std_logic_vector(CFG_NRVEX-1 downto 0);
  signal rctrl2any_traceStall     : std_logic;
  
  -- Misc.
  signal dipsw_int                : std_logic_vector(7 downto 0);
  
begin
  
  ------------------------------------------------------------------------------
  -- Clocking stuff
  ------------------------------------------------------------------------------
  
  -- 125 MHz clock from the Ethernet oscillator.
  gtxclk0 : entity work.gtxclk
    port map (
      clk_p   => gmiiclk_p,
      clk_n   => gmiiclk_n,
      clkint  => clk125,
      clkout  => open
    );
  
  -- 33 MHz clock from the system ACE oscillator.
  clk_33_pad : clkpad
    generic map (
      level   => cmos,
      voltage => x25v,
      tech    => padtech
    )
    port map (
      pad     => clk_33,
      o       => clk33
    );
  
  -- PLL lock signal.
  lock <= phy_init_done;
  led(1) <= phy_init_done;
  
  
  ------------------------------------------------------------------------------
  -- Reset stuff
  ------------------------------------------------------------------------------
  
  reset_block: block is

    signal lockTimeoutRst   : std_logic;
    signal lockTimeoutA     : unsigned(12 downto 0) := (others => '0');
    signal lockTimeoutB     : unsigned(13 downto 0) := (others => '0');
    signal lockTimeout      : std_logic;
    signal resetOrTimeout   : std_logic;

    -- lockTimeoutRst and lockTimeout cross two independent clock domains.
    -- Their timing is completely irrelevant because they're treated as
    -- asynchronous signals, so we need to disable timing checking for these
    -- signals. To do that, we can't have them be optimized away, so we need
    -- to attach the KEEP property to them. The actual TIG constraint has to
    -- be placed in the UCF file.
    attribute KEEP                    : string;
    attribute KEEP of lockTimeoutRst  : signal is "TRUE";
    attribute KEEP of lockTimeout     : signal is "TRUE";

  begin

    -- Generate reset signal for the clock lock/PHY init timeout.
    lockTimeoutRst <= reset or lock;

    -- Generate the lock/PHY timeout counters. Use the clkace 33 MHz clock
    -- signal for this instead of clkm, because clkace always runs,
    -- whereas clkm comes from an MMCM in the MIG, which is reset when
    -- we generate a timeout.
    lock_timeout_proc: process (clk33) is
    begin
      if rising_edge(clk33) then
        if lockTimeoutRst = '1' then
          lockTimeoutA  <= (others => '0');
          lockTimeoutB  <= (others => '0');
          lockTimeout   <= '0';
        else
          if lockTimeoutA(12) = '0' then
            lockTimeoutA <= lockTimeoutA + 1;
          else
            lockTimeoutA <= (others => '0');
            if lockTimeoutB(13) = '0' then
              lockTimeoutB <= lockTimeoutB + 1;
            else
              lockTimeoutB <= (others => '0');
            end if;
          end if;
          lockTimeout <= lockTimeoutB(12) and lockTimeoutB(11)
                     and lockTimeoutB(10) and lockTimeoutB(9);
        end if;
      end if;
    end process;

    -- Combine the incoming reset signal with the lock timeout.
    resetOrTimeout <= reset or lockTimeout;

    -- Original reset generator.
    rst0 : rstgen
      generic map (
        acthigh   => 1
      )
      port map (
        rstin     => resetOrTimeout,
        clk       => clkm,
        clklock   => lock,
        rstout    => rstn,
        rstoutraw => rstraw
      );

  end block;
  
  
  ------------------------------------------------------------------------------
  -- Bus control
  ------------------------------------------------------------------------------
  -- Masters:
  --   0: r-VEX lane group 0
  --   1: r-VEX lane group 1
  --   2: r-VEX lane group 2
  --   3: r-VEX lane group 3
  --   4: ahbjtag
  --   5: bus2ahb (debug UART)
  --
  -- AHB slaves:
  --   0: ahb2mig     0x00000000..0x3FFFFFFF
  --   1: apbctrl     0x80000000..0x8FFFFFFF
  --   2: ahb2bus     0xD0000000..0xDFFFFFFF
  --
  -- APB slaves:
  --   0: gpio        0x80000500..0x800005FF
  --
  -- r-VEX bus slaves:
  --   r-VEX i        0xD00i0000..0xD00iFFFF
  --   debug UART     0xD1000000..0xD1000007                IRQ 2
  --   irq controller 0xD2000000..0xD20007FF
  --
  -- Memory map:
  --    .-----------.---------------.------------.-----.----------------------------------------------.
  --    | Periph.   | Address space | Bw. compat.| IRQ | Description                                  |
  --    |- - - - - -+- - - - - - - - `------. - -+- - -+- - - - - - - - - - - - - - - - - - - - - - - |
  --    | ahbmig    | 0x00000000..0x3FFFFFFF | * |     | Main memory                                  |
  --    | ---       | 0x40000000..0x800004FF |   |     | ---                                          |
  --    | gpio      | 0x80000500..0x800005FF |   |     | Switches, buttons, LEDs                      |
  --    | ---       | 0x80000600..0xCFFFFFFF |   |     | ---                                          |
  --    | rvex      | 0xD0000000..0xD0001FFF | * |     | Primary r-VEX core                           |
  --    | trace     | 0xD0002000..0xD0003FFF | * |     | Trace buffer for primary r-VEX core          |
  --    | ---       | 0xD0004000..0xD00FFFFF |   |     | ---                                          |
  --    | rvex      | 0xD0100000..0xD0101FFF | * |     | Second r-VEX core (if instantiated)          |
  --    | trace     | 0xD0102000..0xD0103FFF | * |     | Trace buffer for second r-VEX core           |
  --    | ---       | 0xD0104000..0xD01FFFFF |   |     | ---                                          |
  --    | ...       | ...................... |   |     | ...                                          |
  --    | ---       | 0xD0x04000..0xD0FFFFFF |   |     | ---                                          |
  --    | dbguart   | 0xD1000000..0xD1000007 | * | 2   | Debug UART                                   |
  --    | ---       | 0xD1000008..0xD1FFFFFF |   |     | ---                                          |
  --    | irq ctrl  | 0xD2000000..0xD20007FF |   | 1   | Interrupt controller and timer               |
  --    | ---       | 0xD2000800..0xD2FFFFFF |   |     | ---                                          |
  --    | busy_cnt  | 0xD3000000..0xD3000003 |   |     | Overall cycle counter                        |
  --    | ---       | 0xD3000004..0xFFFFFFFF |   |     | ---                                          |
  --    '-----------'------------------------'---'-----'----------------------------------------------'
  --
  -- Bw. compat.: backwards compatible with old grlib platform.
  
  -- AHB controller.
  ahb : ahbctrl
    generic map (
      rrobin                    => 1,
      nahbm                     => CFG_NLG+2,
      nahbs                     => 3
    )
    port map (
      rst                       => rstn,
      clk                       => clkm,
      msti                      => ahbmi,
      msto                      => ahbmo,
      slvi                      => ahbsi,
      slvo                      => ahbso
    );
  
  -- APB bridge.
  apb : apbctrl
    generic map (
      hindex                    => 1,
      haddr                     => 16#800#,
      hmask                     => 16#F00#,
      nslaves                   => 1
    )
    port map (
      rst                       => rstn,
      clk                       => clkm,
      ahbi                      => ahbsi,
      ahbo                      => ahbso(1),
      apbi                      => apbi,
      apbo                      => apbo
    );
  
  
  -- r-VEX bus bridge.
  rvex_bus_bridge_block: block is

    signal reset        : std_logic;
    signal clk          : std_logic;
    
    -- Busses between the demuxer and the bus stages.
    signal rvbsi_s      : bus_mst2slv_array(0 to N_RVB_SLAVES - 1);
    signal rvbso_s      : bus_slv2mst_array(0 to N_RVB_SLAVES - 1);
  
    function addr_map return addrRangeAndMapping_array is
      variable retval : addrRangeAndMapping_array(0 to N_RVB_SLAVES - 1);
      variable i : natural;
    begin
      i := 0;
      
      -- Processors.
      for c in 0 to CFG_NRVEX - 1 loop
        retval(i) := addrRangeAndMap(
          match => "------00" & std_logic_vector(to_unsigned(c, 4)) & "----" & "--------" & "--------"
        );
        i := i + 1;
      end loop;
      
      -- Debug UART.
      retval(i) := addrRangeAndMap(
        match => "------01" & "--------" & "--------" & "--------"
      );
      i := i + 1;
      
      -- Interrupt controller/timer.
      retval(i) := addrRangeAndMap(
        match => "------10" & "--------" & "--------" & "--------"
      );
      i := i + 1;
      
      -- Busy LED/performance counter.
      retval(i) := addrRangeAndMap(
        match => "------11" & "--------" & "--------" & "--------"
      );
      i := i + 1;
      
      return retval;
    end function;

  begin

    reset <= not rstn;
    clk <= clkm;

    -- Instantiate the bus bridge.
    rvex_bus_bridge_inst: entity rvex.ahb2bus
      generic map (
        AHB_INDEX       => 2,
        AHB_ADDR        => 16#D00#,
        AHB_MASK        => 16#F00#,
        AHB_VENDOR_ID   => VENDOR_TUDELFT,
        AHB_DEVICE_ID   => TUDELFT_BRIDGE
      )
      port map (
        reset           => reset,
        clk             => clk,
        ahb2bridge      => ahbsi,
        bridge2ahb      => ahbso(2),
        bridge2bus      => rvbmo,
        bus2bridge      => rvbmi
      );

    -- Instantiate the demuxer.
    rvex_bus_bridge_demux: entity rvex.bus_demux
      generic map (
        ADDRESS_MAP     => addr_map
      )
      port map (
        reset           => reset,
        clk             => clk,
        clkEn           => '1',
        mst2demux       => rvbmo,
        demux2mst       => rvbmi,
        demux2slv       => rvbsi_s,
        slv2demux       => rvbso_s
      );
    
    -- Generate the bus stage registers to make routing a bit easier.
    rvex_bus_stages: for i in 0 to N_RVB_SLAVES - 1 generate
      rvex_bus_stage: entity rvex.bus_stage
        port map (
          reset           => reset,
          clk             => clk,
          clkEn           => '1',
          mst2stage       => rvbsi_s(i),
          stage2mst       => rvbso_s(i),
          stage2slv       => rvbsi(i),
          slv2stage       => rvbso(i)
        );
    end generate;
    
  end block;
  
  
  ------------------------------------------------------------------------------
  -- r-VEX processor
  ------------------------------------------------------------------------------
  
  rvsys_gen: for i in 0 to CFG_NRVEX-1 generate
    
    -- Calculate the lIND of the current core depending on the number of
    -- lane groups of all previous cores.
    function CALC_LIND return integer is
      variable LIND : integer := 0;
    begin
      for index in 0 to i-1 loop
        LIND := LIND + 2**CFG_RVEX_CFG(index).core.numLaneGroupsLog2;
      end loop;
      return LIND;
    end function;
    
    -- Calculate the CIND of the current core depending on the number of
    -- contexts of all previous cores.
    function CALC_CIND return integer is
      variable CIND : integer := 0;
    begin
      for index in 0 to i-1 loop
        CIND := CIND + 2**CFG_RVEX_CFG(index).core.numContextsLog2;
      end loop;
      return CIND;
    end function;
    
    constant LIND : integer := CALC_LIND;
    constant LNUM : integer := 2**CFG_RVEX_CFG(i).core.numLaneGroupsLog2;
    constant CIND : integer := CALC_CIND;
    constant CNUM : integer := 2**CFG_RVEX_CFG(i).core.numContextsLog2;
  begin

    rvsys_inst: entity rvex.rvsys_grlib_rctrl
      generic map (
        CFG                     => CFG_RVEX_CFG(i),
        PLATFORM_TAG            => RVEX_PLATFORM_TAG,
        AHB_MASTER_INDEX_START  => LIND,
        CHECK_MEM               => false,
        CHECK_MEM_FILE          => "ram.srec"
      )
      port map (
        clki                    => clkm,
        rstn                    => rstn,
        ahbmi                   => ahbmi,
        ahbmo                   => ahbmo(LIND+LNUM-1 downto LIND),
        ahbsi                   => ahbsi,
        bus2dgb                 => rvbsi(i),
        dbg2bus                 => rvbso(i),
        rctrl2rv_irq            => irq2rv_irq(CIND+CNUM-1 downto CIND),
        rctrl2rv_irqID          => irq2rv_irqID(CIND+CNUM-1 downto CIND),
        rv2rctrl_irqAck         => rv2irq_irqAck(CIND+CNUM-1 downto CIND),
        rctrl2rv_run            => busy2rv_run(CIND+CNUM-1 downto CIND),
        rv2rctrl_idle           => rv2irq_idle(CIND+CNUM-1 downto CIND),
        rv2rctrl_break          => rv2irq_break(CIND+CNUM-1 downto CIND),
        rv2rctrl_traceStall     => rv2rctrl_traceStall(i),
        rctrl2rv_traceStall     => rctrl2any_traceStall,
        rctrl2rv_reset          => irq2rv_reset(CIND+CNUM-1 downto CIND),
        --rctrl2rv_resetVect      => irq2rv_resetVect(CIND+CNUM-1 downto CIND), -- Use the CFG reset vectors
        rv2rctrl_done           => rv2irq_done(CIND+CNUM-1 downto CIND),
        gpio_dip                => dipsw_int
      );

  end generate;
  
  -- Merge the trace stall signals.
  trace_merge: process (rv2rctrl_traceStall) is
    variable flag : std_logic;
  begin
    flag := '0';
    for i in rv2rctrl_traceStall'range loop
      flag := flag or rv2rctrl_traceStall(i);
    end loop;
    rctrl2any_traceStall <= flag;
  end process;
  
  
  ------------------------------------------------------------------------------
  -- Interrupt controller
  ------------------------------------------------------------------------------
  
  irqctrl_block: block is
    signal reset        : std_logic;
    signal clk          : std_logic;
  begin
    
    reset <= not rstn;
    clk <= clkm;

    irqctrl: entity rvex.periph_irq
      generic map (
        BASE_ADDRESS            => X"D2000000",
        NUM_CONTEXTS            => CFG_NCTXT,
        NUM_IRQ                 => NIRQ,
        CONFIG_PRIO_ENABLE      => 1,
        NESTING_ENABLE          => 1,
        BREAKPOINT_BROADCASTING => 1,
        CONFIG_RVECT_ENABLE     => 1,
        OUTPUT_REGISTER         => 1
      )
      port map (
        
        -- System control.
        reset                   => reset,
        clk                     => clk,
        clkEn                   => '1',
        
        -- r-VEX interface.
        irq2rv_irq              => irq2rv_irq,
        irq2rv_irqID            => irq2rv_irqID,
        rv2irq_irqAck           => rv2irq_irqAck,
        irq2rv_run              => irq2busy_run,
        rv2irq_idle             => rv2irq_idle,
        rv2irq_break            => rv2irq_break,
        rv2irq_traceStall       => rctrl2any_traceStall,
        irq2rv_reset            => irq2rv_reset,
        irq2rv_resetVect        => irq2rv_resetVect,
        rv2irq_done             => rv2irq_done,
       
        -- Interrupt inputs.
        periph2irq              => irq,
        
        -- Bus interface.
        bus2irq                 => rvbsi(CFG_NRVEX+1),
        irq2bus                 => rvbso(CFG_NRVEX+1)
        
      );
    
  end block;
  
  
  ------------------------------------------------------------------------------
  -- Busy LED and total cycle counter
  ------------------------------------------------------------------------------
  
  busy_counter: block is
    signal reset        : std_logic;
    signal clk          : std_logic;
    signal idle_counter : std_logic_vector(6 downto 0);
    signal busy         : std_logic;
    signal perf_counter : rvex_data_type;
    signal run          : std_logic;
  begin
    
    reset <= not rstn;
    clk <= clkm;
    
    reg_proc: process (clk) is
      variable idle : std_logic;
    begin
      if rising_edge(clk) then
        rvbso(CFG_NRVEX+2) <= BUS_SLV2MST_IDLE;
        if reset = '1' then
          idle_counter <= (others => '1');
          busy <= '0';
          perf_counter <= (others => '0');
          run <= '1';
        else
          
          -- Determine whether all cores are idle.
          idle := '1';
          for i in rv2irq_idle'range loop
            idle := idle and rv2irq_idle(i);
          end loop;
          
          -- If all cores are idle, increment the idle counter. If the idle
          -- counter is at max, the system is idle. If one of the cores is not
          -- idle, the system is busy and the idle counter is reset to zero.
          if idle = '0' then
            idle_counter <= (others => '0');
            busy <= '1';
          elsif idle_counter /= "1111111" then
            idle_counter <= std_logic_vector(unsigned(idle_counter) + 1);
            busy <= '1';
          else
            busy <= '0';
          end if;
          
          -- If the system is busy, increment the performance counter.
          if busy = '1' then
            perf_counter <= std_logic_vector(unsigned(perf_counter) + 1);
          end if;
          
          -- Handle reads of the performance counter.
          if rvbsi(CFG_NRVEX+2).readEnable = '1' then
            rvbso(CFG_NRVEX+2).readData <= perf_counter;
            rvbso(CFG_NRVEX+2).ack <= '1';
          end if;
          
          -- Reset the performance counter and the cores if a write occurs,
          -- and write bit 0 to the run flag. If the run flag is cleared, all
          -- cores are artificially paused. This can be used to pause the cores
          -- during program upload and initialization, such that all cores can
          -- be started simultaneously with a single register access.
          if rvbsi(CFG_NRVEX+2).writeEnable = '1' then
            run <= rvbsi(CFG_NRVEX+2).writeData(0);
            perf_counter <= (others => '0');
            rvbso(CFG_NRVEX+2).ack <= '1';
          end if;
          
        end if;
      end if;
    end process;
    
    -- Halt all the cores if the run flag is cleared.
    run_proc: process (irq2busy_run, run) is
    begin
      for i in irq2busy_run'range loop
        busy2rv_run(i) <= irq2busy_run(i) and run;
      end loop;
    end process;
    
    -- Connect LED 7 to the busy signal.
    led(7) <= busy;
    
    -- pragma translate_off
    sim_proc: process is
    begin
      wait until busy = '1';
      wait until busy = '0';
      wait for 100 us;
      assert false report "Simulation complete. It took " & integer'image(to_integer(unsigned(perf_counter))) & " cycles." severity failure;
    end process;
    -- pragma translate_on
    
  end block;
  
  ------------------------------------------------------------------------------
  -- Memory controller
  ------------------------------------------------------------------------------
  -- pragma translate_off
  mig_gen: if not DISABLE_DDR_SIM generate
  begin
  -- pragma translate_on
    
    -- MIG instantiation.
    ddr3ctrl: entity work.mig_37
      generic map (
        SIM_BYPASS_INIT_CAL       => SIM_BYPASS_INIT_CAL,
        CLKOUT_DIVIDE4            => work.config.CFG_MIG_CLK4
      )
      port map (
        clk_ref_p                 => clk_ref_p,
        clk_ref_n                 => clk_ref_n,
        ddr3_dq                   => ddr3_dq,
        ddr3_addr                 => ddr3_addr,
        ddr3_ba                   => ddr3_ba,
        ddr3_ras_n                => ddr3_ras_n,
        ddr3_cas_n                => ddr3_cas_n,
        ddr3_we_n                 => ddr3_we_n,
        ddr3_reset_n              => ddr3_reset_n,
        ddr3_cs_n                 => ddr3_cs_n,
        ddr3_odt                  => ddr3_odt,
        ddr3_cke                  => ddr3_cke,
        ddr3_dm                   => ddr3_dm,
        ddr3_dqs_p                => ddr3_dqs_p,
        ddr3_dqs_n                => ddr3_dqs_n,
        ddr3_ck_p                 => ddr3_ck_p,
        ddr3_ck_n                 => ddr3_ck_n,
        app_wdf_wren              => migi.app_wdf_wren,
        app_wdf_data              => migi.app_wdf_data,
        app_wdf_mask              => migi.app_wdf_mask,
        app_wdf_end               => migi.app_wdf_end,
        app_addr                  => migi.app_addr,
        app_cmd                   => migi.app_cmd,
        app_en                    => migi.app_en,
        app_rdy                   => migo.app_rdy,
        app_wdf_rdy               => migo.app_wdf_rdy,
        app_rd_data               => migo.app_rd_data,
        app_rd_data_valid         => migo.app_rd_data_valid,
        tb_rst                    => open,
        tb_clk                    => clkddr,
        clk_ahb                   => clkm,
        clk100                    => clk100,
        phy_init_done             => phy_init_done,
        sys_rst_13                => reset,
        sys_rst_14                => rstraw
      );
    
    ahb2mig0 : ahb2mig_ml605
      generic map (
        hindex                    => 0,
        haddr                     => 16#000#,
        hmask                     => 16#C00#,
        MHz                       => 400,  -- Only used for sim debug messages.
        Mbyte                     => 1024, -- Only used for sim debug messages.
        nosync                    => boolean'pos(CFG_MIG_CLK4=12) --CFG_CLKDIV/12)
      ) 
      port map (
        rst                       => rstn,
        clk_ahb                   => clkm,
        clk_ddr                   => clkddr,
        ahbsi                     => ahbsi,
        ahbso                     => ahbso(0),
        migi                      => migi,
        migo                      => migo
      );
    
  -- pragma translate_off
  end generate;
  sim_mem_gen: if DISABLE_DDR_SIM generate
    signal reset        : std_logic;
    signal bridge2model : bus_mst2slv_type;
    signal model2bridge : bus_slv2mst_type;
  begin
    reset <= not rstn;
    
    -- Generate 400 MHz clock.
    process is
    begin
      clkddr <= '1';
      wait for 1250 ps;
      clkddr <= '0';
      wait for 1250 ps;
    end process;
    
    -- Generate 100 MHz clock.
    process is
    begin
      clk100 <= '1';
      wait for 5000 ps;
      clk100 <= '0';
      wait for 5000 ps;
    end process;
    
    -- Generate configurable clock (1200 MHz / CFG_MIG_CLK4).
    process is
    begin
      clkm <= '1';
      wait for CFG_MIG_CLK4 * 417 ps;
      clkm <= '0';
      wait for CFG_MIG_CLK4 * 417 ps;
      clkm <= '1';
      wait for CFG_MIG_CLK4 * 416 ps;
      clkm <= '0';
      wait for CFG_MIG_CLK4 * 417 ps;
      clkm <= '1';
      wait for CFG_MIG_CLK4 * 417 ps;
      clkm <= '0';
      wait for CFG_MIG_CLK4 * 416 ps;
    end process;
    
    -- Generate PHY done signal.
    process is
    begin
      phy_init_done <= '0';
      wait for 1 us;
      phy_init_done <= '1';
      wait;
    end process;
    
    -- Connect the DDR simulation model to nothing.
    ddr3_dq      <= (others => 'Z');
    ddr3_dm      <= (others => '0');
    ddr3_addr    <= (others => '0');
    ddr3_ba      <= (others => '0');
    ddr3_ras_n   <= '1';
    ddr3_cas_n   <= '1';
    ddr3_we_n    <= '1';
    ddr3_reset_n <= '0';
    ddr3_cs_n    <= (others => '1');
    ddr3_odt     <= (others => '0');
    ddr3_cke     <= (others => '0');
    ddr3_dqs_p   <= (others => 'Z');
    ddr3_dqs_n   <= (others => 'Z');
    ddr3_ck_p    <= (others => '0');
    ddr3_ck_n    <= (others => '1');
    
    -- Convert the AHB bus slave interface to r-VEX bus.
    mem_bridge_inst: entity rvex.ahb2bus
      generic map (
        AHB_INDEX       => 0,
        AHB_ADDR        => 16#000#,
        AHB_MASK        => 16#C00#,
        AHB_VENDOR_ID   => VENDOR_TUDELFT,
        AHB_DEVICE_ID   => TUDELFT_BRIDGE
      )
      port map (
        reset           => reset,
        clk             => clkm,
        ahb2bridge      => ahbsi,
        bridge2ahb      => ahbso(0),
        bridge2bus      => bridge2model,
        bus2bridge      => model2bridge
      );
    
    -- Simulate the memory.
    mem_model: process is
      variable mem      : rvmem_memoryState_type;
      variable readData : rvex_data_type;
      variable l        : std.textio.line;
      variable c        : character;
    begin
      
      -- Load the srec file into the memory.
      rvmem_clear(mem, '0');
      rvmem_loadSRec(mem, "ram.srec");
      
      -- Initialize the bus output.
      model2bridge <= BUS_SLV2MST_IDLE;
      
      -- Handle memory requests.
      loop
        
        -- Wait for the next clock.
        wait until rising_edge(clkm);
        
        -- If we have a request, delay for some amount of cycles.
        if bridge2model.readEnable = '1' or bridge2model.writeEnable = '1' then
          model2bridge <= BUS_SLV2MST_IDLE;
          model2bridge.busy <= '1';
          wait until rising_edge(clkm);
          wait until rising_edge(clkm);
          wait until rising_edge(clkm);
          wait until rising_edge(clkm);
          wait until rising_edge(clkm);
        end if;
        
        -- Handle the bus request.
        model2bridge <= BUS_SLV2MST_IDLE;
        if bridge2model.readEnable = '1' then
          rvmem_read(mem, bridge2model.address, readData);
          model2bridge.readData <= readData;
          model2bridge.ack <= '1';
        elsif bridge2model.writeEnable = '1' then
          rvmem_write(mem, bridge2model.address, bridge2model.writeData, bridge2model.writeMask);
          model2bridge.ack <= '1';
        end if;
        
      end loop;
      
    end process;
    
  end generate;
  -- pragma translate_on
  ------------------------------------------------------------------------------
  -- GRMON JTAG interface
  ------------------------------------------------------------------------------
  
  ahbjtag_inst: ahbjtag
    generic map (
      tech                      => fabtech,
      hindex                    => CFG_NLG
    )
    port map(
      rst                       => rstn,
      clk                       => clkm,
      tck                       => '0',
      tms                       => '0',
      tdi                       => '0',
      tdo                       => open,
      ahbi                      => ahbmi,
      ahbo                      => ahbmo(CFG_NLG),
      tapo_tck                  => open,
      tapo_tdi                  => open,
      tapo_inst                 => open,
      tapo_rst                  => open,
      tapo_capt                 => open,
      tapo_shft                 => open,
      tapo_upd                  => open,
      tapi_tdo                  => '0',
      trst                      => '1',
      tdoen                     => open,
      tckn                      => '0',
      tapo_tckn                 => open,
      tapo_ninst                => open,
      tapo_iupd                 => open
    );

  
  ------------------------------------------------------------------------------
  -- Debug UART
  ------------------------------------------------------------------------------
  
  -- Debug UART
  rvuartgen : block
    signal reset        : std_logic;
    signal clk          : std_logic;
    signal rx           : std_logic;
    signal tx           : std_logic;
    signal uart2dbg_bus : bus_mst2slv_type;
    signal dbg2uart_bus : bus_slv2mst_type;
  begin

    reset <= not rstn;
    clk <= clkm;

    -- Instantiate the AHB master for the debug UART.
    rvex_uart_mst_inst: entity rvex.bus2ahb
      generic map (
        AHB_MASTER_INDEX  => CFG_NLG + 1,
        AHB_VENDOR_ID     => VENDOR_TUDELFT,
        AHB_DEVICE_ID     => TUDELFT_UART,
        BUS_ERROR_CODE    => X"00000010",
        REQ_ERROR_CODE    => X"00000011"
      )
      port map (
        reset             => reset,
        clk               => clk,
        bus2bridge        => uart2dbg_bus,
        bridge2bus        => dbg2uart_bus,
        bridge2ahb        => ahbmo(CFG_NLG + 1),
        ahb2bridge        => ahbmi
      );

    -- Instantiate the UART.
    rvex_uart_inst: entity rvex.periph_uart
      generic map (
        F_CLK             => real(CLKM_FREQ) * 1000.0,
        F_BAUD            => 115200.0
      )
      port map (
        reset             => reset,
        clk               => clk,
        clkEn             => '1',
        rx                => rx,
        tx                => tx,
        bus2uart          => rvbsi(CFG_NRVEX),
        uart2bus          => rvbso(CFG_NRVEX),
        irq               => irq(2),
        uart2dbg_bus      => uart2dbg_bus,
        dbg2uart_bus      => dbg2uart_bus
      );

    dsurx_pad : inpad generic map (level => cmos, voltage => x25v, tech  => padtech)
      port map (dsurx, rx);
    dsutx_pad : outpad generic map (level => cmos, voltage => x25v, tech => padtech)
      port map (dsutx, tx);
  
    led(2) <= (not rx) or (not tx);
    
  end block;
  
  
  ------------------------------------------------------------------------------
  -- GPIO (LEDs, switches, buttons)
  ------------------------------------------------------------------------------
  
  gpio_block: block is
    signal gpioi                : gpio_in_type;
    signal gpioo                : gpio_out_type;
  begin
    
    gpio_inst: grgpio
      generic map (
        pindex                  => 0,
        paddr                   => 16#005#,
        pmask                   => 16#00F#,
        imask                   => 16#1FFF0000#,
        nbits                   => 29,
        irqgen                  => 0
      )
      port map (
        rst                     => rstn,
        clk                     => clkm,
        apbi                    => apbi,
        apbo                    => apbo(0),
        gpioi                   => gpioi,
        gpioo                   => gpioo
      );
    
    led_pads_1 : outpadv generic map (width => 4, level => cmos, voltage => x25v, tech => padtech)
      port map (led(6 downto 3), gpioo.dout(6 downto 3));
    
    led_pads_2 : outpadv generic map (width => 5, level => cmos, voltage => x25v, tech => padtech)
      port map (led(12 downto 8), gpioo.dout(12 downto 8));
    
    dipsw_pad : inpadv generic map (width => 8, level => cmos, voltage => x15v, tech => padtech)
      port map (dipsw, dipsw_int);
    gpioi.din(23 downto 16) <= dipsw_int;
    
    pbtn_pad : inpadv generic map (width => 5, level => cmos, voltage => x15v, tech => padtech)
      port map (pbtn, gpioi.din(28 downto 24));
    
    gpioi.din(1 downto 0) <= "00";
    gpioi.din(15 downto 13) <= "000";
    
  end block;
  
  
end rtl;
