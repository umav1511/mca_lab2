../config.vhd